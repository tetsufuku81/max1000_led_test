-------------------------------------------------------------------------------
-- Project   : MAX1000
-- File      : max1000_led.vhd
-- Title     : MAX1000 Lチカ
--------------------------------------------------------------------------------
--+-----+-----------+-----------------------------------------------------------
-- Ver   Date        Description
--+-----+-----------+-----------------------------------------------------------
-- 00.00 2019/06/23  Created
--+-----+-----------+-----------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;


entity max1000_led is
  port(
    CLK         : in  std_logic;
    LED_o       : out std_logic_vector(7 downto 0)
  );
END max1000_led;


architecture rtl of max1000_led is

--*************************************************************************************************
-- 変数宣言
--*************************************************************************************************
signal  counter                     : std_logic_vector(20 downto 0)     := (others => '0');
signal  led_status                  : std_logic_vector( 7 downto 0)     := "01111111";

begin
---------------------------------------------------------------------------------------------------
-- カウンタ (12MHzで0.1sをカウント)
---------------------------------------------------------------------------------------------------
process(CLK)
begin
  if (CLK'event and CLK = '1') then
    if (counter = "100100100111110000000") then
      counter <= (others => '0');
    else
      counter <= counter + 1;
    end if;

  end if;
end process;

---------------------------------------------------------------------------------------------------
-- LED制御
---------------------------------------------------------------------------------------------------
process(CLK)
begin
  if (CLK'event and CLK = '1') then
    if (counter = "100100100111110000000") then
      led_status <= led_status(6 downto 0) & led_status(7);
    end if;
  end if;
end process;

---------------------------------------------------------------------------------------------------
-- 出力FF
---------------------------------------------------------------------------------------------------
process(CLK)
begin
  if (CLK'event and CLK = '1') then
    LED_o <= led_status;
  end if;
end process;

end rtl;
